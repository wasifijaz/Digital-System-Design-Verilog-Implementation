`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:11:07 03/25/2021
// Design Name:   MUX_4x1
// Module Name:   D:/Education/Semester 6/DSD Lab/Lab 2/Lab2/MUX_4x1_tb.v
// Project Name:  Lab2
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: MUX_4x1
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module MUX_4x1_tb;

	// Inputs
	reg i0;
	reg i1;
	reg i2;
	reg i3;
	reg s1;
	reg s0;

	// Outputs
	wire out;

	// Instantiate the Unit Under Test (UUT)
	MUX_4x1 uut (
		.i0(i0), 
		.i1(i1), 
		.i2(i2), 
		.i3(i3), 
		.s1(s1), 
		.s0(s0), 
		.out(out)
	);

	initial begin
		// Initialize Inputs
		//1
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		//2
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//3
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//4
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//5
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//6
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//7
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//8
		s1 = 0;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;
		
		//9
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
		
		//10
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//11
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//12
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//13
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//14
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//15
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//16
		s1 = 0;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;

		//17
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
		
		//18
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//19
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//20
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//21
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//22
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//23
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//24
		s1 = 0;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;
		
		//25
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
		
		//26
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//27
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//28
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//29
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//30
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//31
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//32
		s1 = 0;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;
		
		//33
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
        
		//34
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//35
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//36
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//37
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//38
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//39
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//40
		s1 = 1;
		s0 = 0;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;
		
		//41
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
		
		//42
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//43
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//44
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//45
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//46
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//47
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//48
		s1 = 1;
		s0 = 0;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;

		//49
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
		
		//50
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//51
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//52
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//53
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//54
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//55
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//56
		s1 = 1;
		s0 = 1;
		i0 = 0;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;
		
		//57
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 0;
		#100;
		
		//58
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 0;
		i3 = 1;
		#100;
		
		//59
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 0;
		#100;
		
		//60
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 0;
		i2 = 1;
		i3 = 1;
		#100;
		
		//61
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 0;
		#100;
		
		//62
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 0;
		i3 = 1;
		#100;
		
		//63
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 0;
		#100;
		
		//64
		s1 = 1;
		s0 = 1;
		i0 = 1;
		i1 = 1;
		i2 = 1;
		i3 = 1;
		#100;
	end
      
endmodule

